*** MODEL Descriptions ***

*** NETLIST Description ***
.LIB "tsmc_025um_model.mod" CMOS_MODELS
.include cmos.sub
X1 out in vdd 0 cmos_inverter

cload out 0 10f
Vdd vdd 0 2.5
Vin in 0 0 pulse 0 2.5 0 10p 10p 1n 2n
*** SIMULATION Commands ***
.op
.tran 10p 5n
*** .include tsmc_025um_model.mod  ***
.end

