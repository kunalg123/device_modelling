*** MODEL Descriptions ***

*** NETLIST Description ***

M1 vdd n1 0 0 nmos W=0.375u L=0.25u

R1 in n1 55

Vdd vdd 0 2.5

Vin in 0 2.5

*** SIMULATION Commands ***

.op

.dc Vin 0 2.5 0.1 Vdd 0 2.5 2.5

*** .include mosis_1um_model.mod ***

.LIB "tsmc_025um_model.mod" CMOS_MODELS

.end


